module rotateN_tb;